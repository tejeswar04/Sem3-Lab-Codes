`timescale 1ns/1ns
`include "question2.v"
module question2_tb;
reg x1,x2,x3,x4;
wire f;
question2 q2(x1,x2,x3,x4,f);
initial begin
$dumpfile("question2_tb.vcd");
$dumpvars(0,question2_tb);
	x1=0;
	x2=0;
	x3=0;
	x4=0;
	#5; 
	x1=0;
	x2=0;
	x3=0;
	x4=1;
	#5; 
	x1=0;
	x2=0;
	x3=1;
	x4=0;
	#5; 
	x1=0;
	x2=0;
	x3=1;
	x4=1;
	#5; 
	x1=0;
	x2=1;
	x3=0;
	x4=0;
	#5; 
	x1=0;
	x2=1;
	x3=0;
	x4=1;
	#5; 
	x1=0;
	x2=1;
	x3=1;
	x4=0;
	#5; 
	x1=0;
	x2=1;
	x3=1;
	x4=1;
	#5; 
	x1=1;
	x2=0;
	x3=0;
	x4=0;
	#5; 
	x1=1;
	x2=0;
	x3=0;
	x4=1;
	#5; 
	x1=1;
	x2=0;
	x3=1;
	x4=0;
	#5; 
	x1=1;
	x2=0;
	x3=1;
	x4=1;
	#5; 
	x1=1;
	x2=1;
	x3=0;
	x4=0;
	#5; 
	x1=1;
	x2=1;
	x3=0;
	x4=1;
	#5; 
	x1=1;
	x2=1;
	x3=1;
	x4=0;
	#5; 
	x1=1;
	x2=1;
	x3=1;
	x4=1;
	#5; 
	$display("Completed");
end
endmodule
