`timescale 1ns/1ns
`include "q1a.v"
module q1a_tb;
reg x1,x2,x3,x4;
wire f;
q1a q1a1(x1,x2,x3,x4,f);
initial begin
	$dumpfile("q1a_tb.vcd");
	$dumpvars(0,q1a_tb);
	x1=0;
	x2=0;
	x3=0;
	x4=0;
	#5; 
	x1=0;
	x2=0;
	x3=0;
	x4=1;
	#5; 
	x1=0;
	x2=0;
	x3=1;
	x4=0;
	#5; 
	x1=0;
	x2=0;
	x3=1;
	x4=1;
	#5; 
	x1=0;
	x2=1;
	x3=0;
	x4=0;
	#5; 
	x1=0;
	x2=1;
	x3=0;
	x4=1;
	#5; 
	x1=0;
	x2=1;
	x3=1;
	x4=0;
	#5; 
	x1=0;
	x2=1;
	x3=1;
	x4=1;
	#5; 
	x1=1;
	x2=0;
	x3=0;
	x4=0;
	#5; 
	x1=1;
	x2=0;
	x3=0;
	x4=1;
	#5; 
	x1=1;
	x2=0;
	x3=1;
	x4=0;
	#5; 
	x1=1;
	x2=0;
	x3=1;
	x4=1;
	#5; 
	x1=1;
	x2=1;
	x3=0;
	x4=0;
	#5; 
	x1=1;
	x2=1;
	x3=0;
	x4=1;
	#5; 
	x1=1;
	x2=1;
	x3=1;
	x4=0;
	#5; 
	x1=1;
	x2=1;
	x3=1;
	x4=1;
	#5;
	$display("Test Completed");
end
endmodule
