`timescale 1ns/1ns
`include "Mux16_1.v"
module Mux16_1_tb;
reg [0:15]W;
reg [3:0]S;
wire f;
Mux16_1 M1(W,S,f);
initial begin
$dumpfile("Mux16_1_tb.vcd");
$dumpvars(0,Mux16_1_tb);
	W=16'b1010101010101010;
	S=0;
	#20;
	W=16'b1010101010101010;
	S=1;
	#20;
	W=16'b1010101010101010;
	S=2;
	#20;
	W=16'b1010101010101010;
	S=3;
	#20;
	W=16'b1010101010101010;
	S=4;
	#20;
	W=16'b1010101010101010;
	S=5;
	#20;
	W=16'b1010101010101010;
	S=6;
	#20;
	W=16'b1010101010101010;
	S=7;
	#20;
	W=16'b1010101010101010;
	S=8;
	#20;
	W=16'b1010101010101010;
	S=9;
	#20;
	W=16'b1010101010101010;
	S=10;
	#20;
	W=16'b1010101010101010;
	S=11;
	#20;
	W=16'b1010101010101010;
	S=12;
	#20;
	W=16'b1010101010101010;
	S=13;
	#20;
	W=16'b1010101010101010;
	S=14;
	#20;
	W=16'b1010101010101010;
	S=15;
	#20;
end
endmodule
