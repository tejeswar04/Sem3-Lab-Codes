module add1(x1,x2,x3,f1,f2);
input x1,x2,x3;
output f1,f2;

